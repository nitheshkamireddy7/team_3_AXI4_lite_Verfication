class axi_coverage;

  

endclass
