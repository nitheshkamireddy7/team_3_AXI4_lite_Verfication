class environment;
  virtual axi_if axi;
  function new(axi_if axi);
    this.axi = axi;
  endfunction

  
