class read_generator;
  mailbox #(read_txn) rbox;
  read_txn rtx;
